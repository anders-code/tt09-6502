/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_anders_tt_6502 (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // All output pins must be assigned. If not used, assign to 0.
//  assign uo_out  = ui_in + uio_in;  // Example: ou_out is the sum of ui_in and uio_in
  assign uio_out = 0;
  assign uio_oe  = 0;

  reg [7:0]mem[16];
  reg [7:0]memout;
  always_ff @(posedge clk) begin
      if (ui_in[7])
          mem[ui_in[3:0]] <= uio_in[7:0];
      memout <= mem[ui_in[3:0]];
  end

  assign uo_out = memout;

  // List all unused inputs to prevent warnings
  wire _unused = &{ui_in[6:4], ena, clk, rst_n, 1'b0};

endmodule
